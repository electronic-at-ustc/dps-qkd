----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:21:20 11/26/2014 
-- Design Name: 
-- Module Name:    div16 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- megafunction wizard: %LPM_DIVIDE% 
-- GENERATION: STANDARD 
-- VERSION: WM1.0 
-- MODULE: lpm_divide  
 
-- ============================================================ 
-- File Name: div16.vhd 
-- Megafunction Name(s): 
-- 			lpm_divide 
-- ============================================================ 
-- ************************************************************ 
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE! 
-- 
-- 6.0 Build 178 04/27/2006 SJ Full Version 
-- ************************************************************ 
 
 
--Copyright (C) 1991-2006 Altera Corporation 
--Your use of Altera Corporation's design tools, logic functions  
--and other software and tools, and its AMPP partner logic  
--functions, and any output files any of the foregoing  
--(including device programming or simulation files), and any  
--associated documentation or information are expressly subject  
--to the terms and conditions of the Altera Program License  
--Subscription Agreement, Altera MegaCore Function License  
--Agreement, or other applicable license agreement, including,  
--without limitation, that your use is for the sole purpose of  
--programming logic devices manufactured by Altera and sold by  
--Altera or its authorized distributors.  Please refer to the  
--applicable agreement for further details. 
 
 
LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
 
LIBRARY lpm; 
USE lpm.all; 
 
ENTITY div16 IS 
	PORT 
	( 
		clock		: IN STD_LOGIC ; 
		denom		: IN STD_LOGIC_VECTOR (8 DOWNTO 0); 
		numer		: IN STD_LOGIC_VECTOR (17 DOWNTO 0); 
		quotient		: OUT STD_LOGIC_VECTOR (17 DOWNTO 0); 
		remain		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0) 
	); 
END div16; 
 
 
ARCHITECTURE SYN OF div16 IS 
 
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (17 DOWNTO 0); 
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (8 DOWNTO 0); 
 
 
 
	COMPONENT lpm_divide 
	GENERIC ( 
		lpm_drepresentation		: STRING; 
		lpm_hint		: STRING; 
		lpm_nrepresentation		: STRING; 
		lpm_pipeline		: NATURAL; 
		lpm_type		: STRING; 
		lpm_widthd		: NATURAL; 
		lpm_widthn		: NATURAL 
	); 
	PORT ( 
			denom	: IN STD_LOGIC_VECTOR (8 DOWNTO 0); 
			clock	: IN STD_LOGIC ; 
			quotient	: OUT STD_LOGIC_VECTOR (17 DOWNTO 0); 
			remain	: OUT STD_LOGIC_VECTOR (8 DOWNTO 0); 
			numer	: IN STD_LOGIC_VECTOR (17 DOWNTO 0) 
	); 
	END COMPONENT; 
 
BEGIN 
	quotient    <= sub_wire0(17 DOWNTO 0); 
	remain    <= sub_wire1(8 DOWNTO 0); 
 
	lpm_divide_component : lpm_divide 
	GENERIC MAP ( 
		lpm_drepresentation => "UNSIGNED", 
		lpm_hint => "LPM_REMAINDERPOSITIVE=TRUE", 
		lpm_nrepresentation => "UNSIGNED", 
		lpm_pipeline => 4, 
		lpm_type => "LPM_DIVIDE", 
		lpm_widthd => 9, 
		lpm_widthn => 18 
	) 
	PORT MAP ( 
		denom => denom, 
		clock => clock, 
		numer => numer, 
		quotient => sub_wire0, 
		remain => sub_wire1 
	); 
 
 
 
END SYN; 
 
-- ============================================================ 
-- CNX file retrieval info 
-- ============================================================ 
-- Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE" 
-- Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1" 
-- Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "1" 
-- Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2" 
-- Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED" 
-- Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE" 
-- Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED" 
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "4" 
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE" 
-- Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "9" 
-- Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "18" 
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock 
-- Retrieval info: USED_PORT: denom 0 0 9 0 INPUT NODEFVAL denom[8..0] 
-- Retrieval info: USED_PORT: numer 0 0 18 0 INPUT NODEFVAL numer[17..0] 
-- Retrieval info: USED_PORT: quotient 0 0 18 0 OUTPUT NODEFVAL quotient[17..0] 
-- Retrieval info: USED_PORT: remain 0 0 9 0 OUTPUT NODEFVAL remain[8..0] 
-- Retrieval info: CONNECT: @numer 0 0 18 0 numer 0 0 18 0 
-- Retrieval info: CONNECT: @denom 0 0 9 0 denom 0 0 9 0 
-- Retrieval info: CONNECT: quotient 0 0 18 0 @quotient 0 0 18 0 
-- Retrieval info: CONNECT: remain 0 0 9 0 @remain 0 0 9 0 
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0 
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all 
-- Retrieval info: GEN_FILE: TYPE_NORMAL div16.vhd TRUE 
-- Retrieval info: GEN_FILE: TYPE_NORMAL div16.inc FALSE 
-- Retrieval info: GEN_FILE: TYPE_NORMAL div16.cmp FALSE 
-- Retrieval info: GEN_FILE: TYPE_NORMAL div16.bsf FALSE 
-- Retrieval info: GEN_FILE: TYPE_NORMAL div16_inst.vhd FALSE 
